

/*
Modelo de ALU para el microprocesador de 8 bits.
*/

